`include "includes.sv"

module top;
    
    testbench   tb();

endmodule

 `include "testbench.sv"
 `include "clk_gen.sv"
 `include "approx_2x2.sv"
 `include "approx_4x4.sv"
 `include "precise_2x2.sv"
 `include "precise_4x4.sv"
 `include "approx_8x8.sv"
 `include "approx_16x16.sv"
